module led_top (
    input  logic        clk,
    input  logic        rst,          // Active high
    input  logic [31:0] csr_addr,
    input  logic [31:0] csr_wdata,
    input  logic        csr_write,
    output logic [31:0] csr_rdata,
    output logic        led_out
);

    // Internal signals for the "passthrough" bus
    logic        s_cpuif_req;
    logic        s_cpuif_req_is_wr;
    logic [2:0]  s_cpuif_addr;
    logic [31:0] s_cpuif_wr_data;
    logic [31:0] s_cpuif_wr_biten;
    logic        s_cpuif_rd_ack;
    logic [31:0] s_cpuif_rd_data;

    // Register output structure
    led_regs_pkg::led_regs__out_t hwif_out;

    // Simple adapter: each operation lasts 1 cycle
    assign s_cpuif_req       = csr_write || (csr_addr !== 32'hx);
    assign s_cpuif_req_is_wr = csr_write;
    assign s_cpuif_addr      = csr_addr[4:2];   // Adjust according to address size
    assign s_cpuif_wr_data   = csr_wdata;
    assign s_cpuif_wr_biten  = 32'hFFFF_FFFF;   // Write all bits
    assign csr_rdata         = s_cpuif_rd_data;

    // Instance of the register block generated by PeakRDL
    led_regs regs_inst (
        .clk                  (clk),
        .rst                  (rst),
        .s_cpuif_req          (s_cpuif_req),
        .s_cpuif_req_is_wr    (s_cpuif_req_is_wr),
        .s_cpuif_addr         (s_cpuif_addr),
        .s_cpuif_wr_data      (s_cpuif_wr_data),
        .s_cpuif_wr_biten     (s_cpuif_wr_biten),
        .s_cpuif_req_stall_wr (), // Not used
        .s_cpuif_req_stall_rd (), // Not used
        .s_cpuif_rd_ack       (s_cpuif_rd_ack),
        .s_cpuif_rd_err       (), // Not used
        .s_cpuif_rd_data      (s_cpuif_rd_data),
        .s_cpuif_wr_ack       (), // Not used
        .s_cpuif_wr_err       (), // Not used
        .hwif_out             (hwif_out)
    );

    // Instance of the functional block
    led_controller core_inst (
        .i_clk        (clk),
        .i_rst_n      (~rst),
        .i_enable     (hwif_out.control_inst.ENABLE.value),
        .i_blink_rate (hwif_out.control_inst.BLINK_RATE.value),
        .o_led_out    (led_out)
    );

endmodule
